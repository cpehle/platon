module t1(input logic [31:0] a,
          output logic [31:0] b);
   assign b = a;
endmodule
